//
// t9990_blit_bitmask.sv
//
// BSD 3-Clause License
// 
// Copyright (c) 2024, Shinobu Hashimoto
// 
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
// 
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
// 
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
// 
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
// 
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//

`default_nettype none

/***************************************************************
 * ビットマスク
 ***************************************************************/
module T9990_BLIT_BITMASK (
    input wire          CLK,
    input wire [15:0]   WM,
    input wire [1:0]    CLRM,
    input wire          DIX,
    input wire [3:0]    OFFSET,
    input wire [4:0]    COUNT,
    output reg [31:0]   BIT_MASK
);
    /***************************************************************
     * テーブルから BIT MASK を取得
     ***************************************************************/
    logic [31:0] out_2bpp;
    T9990_BLIT_BITMASK_2BPP u_2bpp (
        .CLK,
        .DIX,
        .OFFSET(OFFSET[3:0]),
        .COUNT(COUNT[4] ? 4'd0 : COUNT[3:0]),
        .OUT(out_2bpp)
    );

    logic [31:0] out_4bpp;
    T9990_BLIT_BITMASK_4BPP u_4bpp (
        .CLK,
        .DIX,
        .OFFSET(OFFSET[2:0]),
        .COUNT(COUNT[4:3] ? 3'd0 : COUNT[2:0]),
        .OUT(out_4bpp)
    );

    logic [31:0] out_8bpp;
    T9990_BLIT_BITMASK_8BPP u_8bpp (
        .CLK,
        .DIX,
        .OFFSET(OFFSET[1:0]),
        .COUNT(COUNT[4:2] ? 2'd0 : COUNT[1:0]),
        .OUT(out_8bpp)
    );

    logic [31:0] out_16bpp;
    T9990_BLIT_BITMASK_16BPP u_16bpp (
        .CLK,
        .DIX,
        .OFFSET(OFFSET[0:0]),
        .COUNT(COUNT[4:1] ? 1'd0 : COUNT[0:0]),
        .OUT(out_16bpp)
    );

    /***************************************************************
     * WM レジスタでマスク
     ***************************************************************/
    always_ff @(posedge CLK) begin
        if(COUNT == 0) begin
            BIT_MASK <= 0;
        end
        else begin
            case (CLRM)
                T9990_REG::CLRM_2BPP:   BIT_MASK <= out_2bpp  & {WM[7:0], WM[15:8], WM[7:0], WM[15:8]};  // ビッグエンディアンで出力するので WM を入れ替え
                T9990_REG::CLRM_4BPP:   BIT_MASK <= out_4bpp  & {WM[7:0], WM[15:8], WM[7:0], WM[15:8]};
                T9990_REG::CLRM_8BPP:   BIT_MASK <= out_8bpp  & {WM[7:0], WM[15:8], WM[7:0], WM[15:8]};
                T9990_REG::CLRM_16BPP:  BIT_MASK <= out_16bpp & {WM[7:0], WM[15:8], WM[7:0], WM[15:8]};
            endcase
        end
    end
endmodule

/***************************************************************
 * 2BPP テーブル
 ***************************************************************/
module T9990_BLIT_BITMASK_2BPP (
    input wire          CLK,
    input wire          DIX,
    input wire [3:0]    OFFSET,
    input wire [3:0]    COUNT,
    output reg [31:0]   OUT
)/* synthesis syn_romstyle="block_rom" */;
    always_ff @(posedge CLK) begin
        case ({DIX,COUNT[3:0],OFFSET[3:0]})
        	9'b0_0001_0000:  	OUT <= 32'b11000000000000000000000000000000;
	        9'b0_0010_0000:  	OUT <= 32'b11110000000000000000000000000000;
    	    9'b0_0011_0000:  	OUT <= 32'b11111100000000000000000000000000;
    	    9'b0_0100_0000:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b0_0101_0000:  	OUT <= 32'b11111111110000000000000000000000;
	        9'b0_0110_0000:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b0_0111_0000:  	OUT <= 32'b11111111111111000000000000000000;
	        9'b0_1000_0000:  	OUT <= 32'b11111111111111110000000000000000;
    	    9'b0_1001_0000:  	OUT <= 32'b11111111111111111100000000000000;
    	    9'b0_1010_0000:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b0_1011_0000:  	OUT <= 32'b11111111111111111111110000000000;
	        9'b0_1100_0000:  	OUT <= 32'b11111111111111111111111100000000;
        	9'b0_1101_0000:  	OUT <= 32'b11111111111111111111111111000000;
	        9'b0_1110_0000:  	OUT <= 32'b11111111111111111111111111110000;
    	    9'b0_1111_0000:  	OUT <= 32'b11111111111111111111111111111100;
    	    9'b0_0000_0000:  	OUT <= 32'b11111111111111111111111111111111;

        	9'b0_0001_0001:  	OUT <= 32'b00110000000000000000000000000000;
	        9'b0_0010_0001:  	OUT <= 32'b00111100000000000000000000000000;
    	    9'b0_0011_0001:  	OUT <= 32'b00111111000000000000000000000000;
    	    9'b0_0100_0001:  	OUT <= 32'b00111111110000000000000000000000;
        	9'b0_0101_0001:  	OUT <= 32'b00111111111100000000000000000000;
	        9'b0_0110_0001:  	OUT <= 32'b00111111111111000000000000000000;
        	9'b0_0111_0001:  	OUT <= 32'b00111111111111110000000000000000;
	        9'b0_1000_0001:  	OUT <= 32'b00111111111111111100000000000000;
    	    9'b0_1001_0001:  	OUT <= 32'b00111111111111111111000000000000;
    	    9'b0_1010_0001:  	OUT <= 32'b00111111111111111111110000000000;
        	9'b0_1011_0001:  	OUT <= 32'b00111111111111111111111100000000;
	        9'b0_1100_0001:  	OUT <= 32'b00111111111111111111111111000000;
        	9'b0_1101_0001:  	OUT <= 32'b00111111111111111111111111110000;
	        9'b0_1110_0001:  	OUT <= 32'b00111111111111111111111111111100;
    	    9'b0_1111_0001:  	OUT <= 32'b00111111111111111111111111111111;
    	    9'b0_0000_0001:  	OUT <= 32'b00111111111111111111111111111111;

        	9'b0_0001_0010:  	OUT <= 32'b00001100000000000000000000000000;
	        9'b0_0010_0010:  	OUT <= 32'b00001111000000000000000000000000;
    	    9'b0_0011_0010:  	OUT <= 32'b00001111110000000000000000000000;
    	    9'b0_0100_0010:  	OUT <= 32'b00001111111100000000000000000000;
        	9'b0_0101_0010:  	OUT <= 32'b00001111111111000000000000000000;
	        9'b0_0110_0010:  	OUT <= 32'b00001111111111110000000000000000;
        	9'b0_0111_0010:  	OUT <= 32'b00001111111111111100000000000000;
	        9'b0_1000_0010:  	OUT <= 32'b00001111111111111111000000000000;
    	    9'b0_1001_0010:  	OUT <= 32'b00001111111111111111110000000000;
    	    9'b0_1010_0010:  	OUT <= 32'b00001111111111111111111100000000;
        	9'b0_1011_0010:  	OUT <= 32'b00001111111111111111111111000000;
	        9'b0_1100_0010:  	OUT <= 32'b00001111111111111111111111110000;
        	9'b0_1101_0010:  	OUT <= 32'b00001111111111111111111111111100;
	        9'b0_1110_0010:  	OUT <= 32'b00001111111111111111111111111111;
    	    9'b0_1111_0010:  	OUT <= 32'b00001111111111111111111111111111;
    	    9'b0_0000_0010:  	OUT <= 32'b00001111111111111111111111111111;

        	9'b0_0001_0011:  	OUT <= 32'b00000011000000000000000000000000;
	        9'b0_0010_0011:  	OUT <= 32'b00000011110000000000000000000000;
    	    9'b0_0011_0011:  	OUT <= 32'b00000011111100000000000000000000;
    	    9'b0_0100_0011:  	OUT <= 32'b00000011111111000000000000000000;
        	9'b0_0101_0011:  	OUT <= 32'b00000011111111110000000000000000;
	        9'b0_0110_0011:  	OUT <= 32'b00000011111111111100000000000000;
        	9'b0_0111_0011:  	OUT <= 32'b00000011111111111111000000000000;
	        9'b0_1000_0011:  	OUT <= 32'b00000011111111111111110000000000;
    	    9'b0_1001_0011:  	OUT <= 32'b00000011111111111111111100000000;
    	    9'b0_1010_0011:  	OUT <= 32'b00000011111111111111111111000000;
        	9'b0_1011_0011:  	OUT <= 32'b00000011111111111111111111110000;
	        9'b0_1100_0011:  	OUT <= 32'b00000011111111111111111111111100;
        	9'b0_1101_0011:  	OUT <= 32'b00000011111111111111111111111111;
	        9'b0_1110_0011:  	OUT <= 32'b00000011111111111111111111111111;
    	    9'b0_1111_0011:  	OUT <= 32'b00000011111111111111111111111111;
    	    9'b0_0000_0011:  	OUT <= 32'b00000011111111111111111111111111;

        	9'b0_0001_0100:  	OUT <= 32'b00000000110000000000000000000000;
	        9'b0_0010_0100:  	OUT <= 32'b00000000111100000000000000000000;
    	    9'b0_0011_0100:  	OUT <= 32'b00000000111111000000000000000000;
    	    9'b0_0100_0100:  	OUT <= 32'b00000000111111110000000000000000;
        	9'b0_0101_0100:  	OUT <= 32'b00000000111111111100000000000000;
	        9'b0_0110_0100:  	OUT <= 32'b00000000111111111111000000000000;
        	9'b0_0111_0100:  	OUT <= 32'b00000000111111111111110000000000;
	        9'b0_1000_0100:  	OUT <= 32'b00000000111111111111111100000000;
    	    9'b0_1001_0100:  	OUT <= 32'b00000000111111111111111111000000;
    	    9'b0_1010_0100:  	OUT <= 32'b00000000111111111111111111110000;
        	9'b0_1011_0100:  	OUT <= 32'b00000000111111111111111111111100;
	        9'b0_1100_0100:  	OUT <= 32'b00000000111111111111111111111111;
        	9'b0_1101_0100:  	OUT <= 32'b00000000111111111111111111111111;
	        9'b0_1110_0100:  	OUT <= 32'b00000000111111111111111111111111;
    	    9'b0_1111_0100:  	OUT <= 32'b00000000111111111111111111111111;
    	    9'b0_0000_0100:  	OUT <= 32'b00000000111111111111111111111111;

        	9'b0_0001_0101:  	OUT <= 32'b00000000001100000000000000000000;
	        9'b0_0010_0101:  	OUT <= 32'b00000000001111000000000000000000;
    	    9'b0_0011_0101:  	OUT <= 32'b00000000001111110000000000000000;
    	    9'b0_0100_0101:  	OUT <= 32'b00000000001111111100000000000000;
        	9'b0_0101_0101:  	OUT <= 32'b00000000001111111111000000000000;
	        9'b0_0110_0101:  	OUT <= 32'b00000000001111111111110000000000;
        	9'b0_0111_0101:  	OUT <= 32'b00000000001111111111111100000000;
	        9'b0_1000_0101:  	OUT <= 32'b00000000001111111111111111000000;
    	    9'b0_1001_0101:  	OUT <= 32'b00000000001111111111111111110000;
    	    9'b0_1010_0101:  	OUT <= 32'b00000000001111111111111111111100;
        	9'b0_1011_0101:  	OUT <= 32'b00000000001111111111111111111111;
	        9'b0_1100_0101:  	OUT <= 32'b00000000001111111111111111111111;
        	9'b0_1101_0101:  	OUT <= 32'b00000000001111111111111111111111;
	        9'b0_1110_0101:  	OUT <= 32'b00000000001111111111111111111111;
    	    9'b0_1111_0101:  	OUT <= 32'b00000000001111111111111111111111;
    	    9'b0_0000_0101:  	OUT <= 32'b00000000001111111111111111111111;

        	9'b0_0001_0110:  	OUT <= 32'b00000000000011000000000000000000;
	        9'b0_0010_0110:  	OUT <= 32'b00000000000011110000000000000000;
    	    9'b0_0011_0110:  	OUT <= 32'b00000000000011111100000000000000;
    	    9'b0_0100_0110:  	OUT <= 32'b00000000000011111111000000000000;
        	9'b0_0101_0110:  	OUT <= 32'b00000000000011111111110000000000;
	        9'b0_0110_0110:  	OUT <= 32'b00000000000011111111111100000000;
        	9'b0_0111_0110:  	OUT <= 32'b00000000000011111111111111000000;
	        9'b0_1000_0110:  	OUT <= 32'b00000000000011111111111111110000;
    	    9'b0_1001_0110:  	OUT <= 32'b00000000000011111111111111111100;
    	    9'b0_1010_0110:  	OUT <= 32'b00000000000011111111111111111111;
        	9'b0_1011_0110:  	OUT <= 32'b00000000000011111111111111111111;
	        9'b0_1100_0110:  	OUT <= 32'b00000000000011111111111111111111;
        	9'b0_1101_0110:  	OUT <= 32'b00000000000011111111111111111111;
	        9'b0_1110_0110:  	OUT <= 32'b00000000000011111111111111111111;
    	    9'b0_1111_0110:  	OUT <= 32'b00000000000011111111111111111111;
    	    9'b0_0000_0110:  	OUT <= 32'b00000000000011111111111111111111;

        	9'b0_0001_0111:  	OUT <= 32'b00000000000000110000000000000000;
	        9'b0_0010_0111:  	OUT <= 32'b00000000000000111100000000000000;
    	    9'b0_0011_0111:  	OUT <= 32'b00000000000000111111000000000000;
    	    9'b0_0100_0111:  	OUT <= 32'b00000000000000111111110000000000;
        	9'b0_0101_0111:  	OUT <= 32'b00000000000000111111111100000000;
	        9'b0_0110_0111:  	OUT <= 32'b00000000000000111111111111000000;
        	9'b0_0111_0111:  	OUT <= 32'b00000000000000111111111111110000;
	        9'b0_1000_0111:  	OUT <= 32'b00000000000000111111111111111100;
    	    9'b0_1001_0111:  	OUT <= 32'b00000000000000111111111111111111;
    	    9'b0_1010_0111:  	OUT <= 32'b00000000000000111111111111111111;
        	9'b0_1011_0111:  	OUT <= 32'b00000000000000111111111111111111;
	        9'b0_1100_0111:  	OUT <= 32'b00000000000000111111111111111111;
        	9'b0_1101_0111:  	OUT <= 32'b00000000000000111111111111111111;
	        9'b0_1110_0111:  	OUT <= 32'b00000000000000111111111111111111;
    	    9'b0_1111_0111:  	OUT <= 32'b00000000000000111111111111111111;
    	    9'b0_0000_0111:  	OUT <= 32'b00000000000000111111111111111111;

        	9'b0_0001_1000:  	OUT <= 32'b00000000000000001100000000000000;
	        9'b0_0010_1000:  	OUT <= 32'b00000000000000001111000000000000;
    	    9'b0_0011_1000:  	OUT <= 32'b00000000000000001111110000000000;
    	    9'b0_0100_1000:  	OUT <= 32'b00000000000000001111111100000000;
        	9'b0_0101_1000:  	OUT <= 32'b00000000000000001111111111000000;
	        9'b0_0110_1000:  	OUT <= 32'b00000000000000001111111111110000;
        	9'b0_0111_1000:  	OUT <= 32'b00000000000000001111111111111100;
	        9'b0_1000_1000:  	OUT <= 32'b00000000000000001111111111111111;
    	    9'b0_1001_1000:  	OUT <= 32'b00000000000000001111111111111111;
    	    9'b0_1010_1000:  	OUT <= 32'b00000000000000001111111111111111;
        	9'b0_1011_1000:  	OUT <= 32'b00000000000000001111111111111111;
	        9'b0_1100_1000:  	OUT <= 32'b00000000000000001111111111111111;
        	9'b0_1101_1000:  	OUT <= 32'b00000000000000001111111111111111;
	        9'b0_1110_1000:  	OUT <= 32'b00000000000000001111111111111111;
    	    9'b0_1111_1000:  	OUT <= 32'b00000000000000001111111111111111;
    	    9'b0_0000_1000:  	OUT <= 32'b00000000000000001111111111111111;

        	9'b0_0001_1001:  	OUT <= 32'b00000000000000000011000000000000;
	        9'b0_0010_1001:  	OUT <= 32'b00000000000000000011110000000000;
    	    9'b0_0011_1001:  	OUT <= 32'b00000000000000000011111100000000;
    	    9'b0_0100_1001:  	OUT <= 32'b00000000000000000011111111000000;
        	9'b0_0101_1001:  	OUT <= 32'b00000000000000000011111111110000;
	        9'b0_0110_1001:  	OUT <= 32'b00000000000000000011111111111100;
        	9'b0_0111_1001:  	OUT <= 32'b00000000000000000011111111111111;
	        9'b0_1000_1001:  	OUT <= 32'b00000000000000000011111111111111;
    	    9'b0_1001_1001:  	OUT <= 32'b00000000000000000011111111111111;
    	    9'b0_1010_1001:  	OUT <= 32'b00000000000000000011111111111111;
        	9'b0_1011_1001:  	OUT <= 32'b00000000000000000011111111111111;
	        9'b0_1100_1001:  	OUT <= 32'b00000000000000000011111111111111;
        	9'b0_1101_1001:  	OUT <= 32'b00000000000000000011111111111111;
	        9'b0_1110_1001:  	OUT <= 32'b00000000000000000011111111111111;
    	    9'b0_1111_1001:  	OUT <= 32'b00000000000000000011111111111111;
    	    9'b0_0000_1001:  	OUT <= 32'b00000000000000000011111111111111;

        	9'b0_0001_1010:  	OUT <= 32'b00000000000000000000110000000000;
	        9'b0_0010_1010:  	OUT <= 32'b00000000000000000000111100000000;
    	    9'b0_0011_1010:  	OUT <= 32'b00000000000000000000111111000000;
    	    9'b0_0100_1010:  	OUT <= 32'b00000000000000000000111111110000;
        	9'b0_0101_1010:  	OUT <= 32'b00000000000000000000111111111100;
	        9'b0_0110_1010:  	OUT <= 32'b00000000000000000000111111111111;
        	9'b0_0111_1010:  	OUT <= 32'b00000000000000000000111111111111;
	        9'b0_1000_1010:  	OUT <= 32'b00000000000000000000111111111111;
    	    9'b0_1001_1010:  	OUT <= 32'b00000000000000000000111111111111;
    	    9'b0_1010_1010:  	OUT <= 32'b00000000000000000000111111111111;
        	9'b0_1011_1010:  	OUT <= 32'b00000000000000000000111111111111;
	        9'b0_1100_1010:  	OUT <= 32'b00000000000000000000111111111111;
        	9'b0_1101_1010:  	OUT <= 32'b00000000000000000000111111111111;
	        9'b0_1110_1010:  	OUT <= 32'b00000000000000000000111111111111;
    	    9'b0_1111_1010:  	OUT <= 32'b00000000000000000000111111111111;
    	    9'b0_0000_1010:  	OUT <= 32'b00000000000000000000111111111111;

        	9'b0_0001_1011:  	OUT <= 32'b00000000000000000000001100000000;
	        9'b0_0010_1011:  	OUT <= 32'b00000000000000000000001111000000;
    	    9'b0_0011_1011:  	OUT <= 32'b00000000000000000000001111110000;
    	    9'b0_0100_1011:  	OUT <= 32'b00000000000000000000001111111100;
        	9'b0_0101_1011:  	OUT <= 32'b00000000000000000000001111111111;
	        9'b0_0110_1011:  	OUT <= 32'b00000000000000000000001111111111;
        	9'b0_0111_1011:  	OUT <= 32'b00000000000000000000001111111111;
	        9'b0_1000_1011:  	OUT <= 32'b00000000000000000000001111111111;
    	    9'b0_1001_1011:  	OUT <= 32'b00000000000000000000001111111111;
    	    9'b0_1010_1011:  	OUT <= 32'b00000000000000000000001111111111;
        	9'b0_1011_1011:  	OUT <= 32'b00000000000000000000001111111111;
	        9'b0_1100_1011:  	OUT <= 32'b00000000000000000000001111111111;
        	9'b0_1101_1011:  	OUT <= 32'b00000000000000000000001111111111;
	        9'b0_1110_1011:  	OUT <= 32'b00000000000000000000001111111111;
    	    9'b0_1111_1011:  	OUT <= 32'b00000000000000000000001111111111;
    	    9'b0_0000_1011:  	OUT <= 32'b00000000000000000000001111111111;

        	9'b0_0001_1100:  	OUT <= 32'b00000000000000000000000011000000;
	        9'b0_0010_1100:  	OUT <= 32'b00000000000000000000000011110000;
    	    9'b0_0011_1100:  	OUT <= 32'b00000000000000000000000011111100;
    	    9'b0_0100_1100:  	OUT <= 32'b00000000000000000000000011111111;
        	9'b0_0101_1100:  	OUT <= 32'b00000000000000000000000011111111;
	        9'b0_0110_1100:  	OUT <= 32'b00000000000000000000000011111111;
        	9'b0_0111_1100:  	OUT <= 32'b00000000000000000000000011111111;
	        9'b0_1000_1100:  	OUT <= 32'b00000000000000000000000011111111;
    	    9'b0_1001_1100:  	OUT <= 32'b00000000000000000000000011111111;
    	    9'b0_1010_1100:  	OUT <= 32'b00000000000000000000000011111111;
        	9'b0_1011_1100:  	OUT <= 32'b00000000000000000000000011111111;
	        9'b0_1100_1100:  	OUT <= 32'b00000000000000000000000011111111;
        	9'b0_1101_1100:  	OUT <= 32'b00000000000000000000000011111111;
	        9'b0_1110_1100:  	OUT <= 32'b00000000000000000000000011111111;
    	    9'b0_1111_1100:  	OUT <= 32'b00000000000000000000000011111111;
    	    9'b0_0000_1100:  	OUT <= 32'b00000000000000000000000011111111;

        	9'b0_0001_1101:  	OUT <= 32'b00000000000000000000000000110000;
	        9'b0_0010_1101:  	OUT <= 32'b00000000000000000000000000111100;
    	    9'b0_0011_1101:  	OUT <= 32'b00000000000000000000000000111111;
    	    9'b0_0100_1101:  	OUT <= 32'b00000000000000000000000000111111;
        	9'b0_0101_1101:  	OUT <= 32'b00000000000000000000000000111111;
	        9'b0_0110_1101:  	OUT <= 32'b00000000000000000000000000111111;
        	9'b0_0111_1101:  	OUT <= 32'b00000000000000000000000000111111;
	        9'b0_1000_1101:  	OUT <= 32'b00000000000000000000000000111111;
    	    9'b0_1001_1101:  	OUT <= 32'b00000000000000000000000000111111;
    	    9'b0_1010_1101:  	OUT <= 32'b00000000000000000000000000111111;
        	9'b0_1011_1101:  	OUT <= 32'b00000000000000000000000000111111;
	        9'b0_1100_1101:  	OUT <= 32'b00000000000000000000000000111111;
        	9'b0_1101_1101:  	OUT <= 32'b00000000000000000000000000111111;
	        9'b0_1110_1101:  	OUT <= 32'b00000000000000000000000000111111;
    	    9'b0_1111_1101:  	OUT <= 32'b00000000000000000000000000111111;
    	    9'b0_0000_1101:  	OUT <= 32'b00000000000000000000000000111111;

        	9'b0_0001_1110:  	OUT <= 32'b00000000000000000000000000001100;
	        9'b0_0010_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_0011_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_0100_1110:  	OUT <= 32'b00000000000000000000000000001111;
        	9'b0_0101_1110:  	OUT <= 32'b00000000000000000000000000001111;
	        9'b0_0110_1110:  	OUT <= 32'b00000000000000000000000000001111;
        	9'b0_0111_1110:  	OUT <= 32'b00000000000000000000000000001111;
	        9'b0_1000_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_1001_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_1010_1110:  	OUT <= 32'b00000000000000000000000000001111;
        	9'b0_1011_1110:  	OUT <= 32'b00000000000000000000000000001111;
	        9'b0_1100_1110:  	OUT <= 32'b00000000000000000000000000001111;
        	9'b0_1101_1110:  	OUT <= 32'b00000000000000000000000000001111;
	        9'b0_1110_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_1111_1110:  	OUT <= 32'b00000000000000000000000000001111;
    	    9'b0_0000_1110:  	OUT <= 32'b00000000000000000000000000001111;

        	9'b0_0001_1111:  	OUT <= 32'b00000000000000000000000000000011;
	        9'b0_0010_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_0011_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_0100_1111:  	OUT <= 32'b00000000000000000000000000000011;
        	9'b0_0101_1111:  	OUT <= 32'b00000000000000000000000000000011;
	        9'b0_0110_1111:  	OUT <= 32'b00000000000000000000000000000011;
        	9'b0_0111_1111:  	OUT <= 32'b00000000000000000000000000000011;
	        9'b0_1000_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_1001_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_1010_1111:  	OUT <= 32'b00000000000000000000000000000011;
        	9'b0_1011_1111:  	OUT <= 32'b00000000000000000000000000000011;
	        9'b0_1100_1111:  	OUT <= 32'b00000000000000000000000000000011;
        	9'b0_1101_1111:  	OUT <= 32'b00000000000000000000000000000011;
	        9'b0_1110_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_1111_1111:  	OUT <= 32'b00000000000000000000000000000011;
    	    9'b0_0000_1111:  	OUT <= 32'b00000000000000000000000000000011;

        	9'b1_0001_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0010_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0011_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0100_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0101_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0110_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0111_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1000_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1001_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1010_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1011_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1100_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1101_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1110_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_1111_0000:  	OUT <= 32'b11000000000000000000000000000000;
        	9'b1_0000_0000:  	OUT <= 32'b11000000000000000000000000000000;

        	9'b1_0001_0001:  	OUT <= 32'b00110000000000000000000000000000;
        	9'b1_0010_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0011_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0100_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0101_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0110_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0111_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1000_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1001_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1010_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1011_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1100_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1101_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1110_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_1111_0001:  	OUT <= 32'b11110000000000000000000000000000;
        	9'b1_0000_0001:  	OUT <= 32'b11110000000000000000000000000000;

        	9'b1_0001_0010:  	OUT <= 32'b00001100000000000000000000000000;
        	9'b1_0010_0010:  	OUT <= 32'b00111100000000000000000000000000;
        	9'b1_0011_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_0100_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_0101_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_0110_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_0111_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1000_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1001_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1010_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1011_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1100_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1101_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1110_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_1111_0010:  	OUT <= 32'b11111100000000000000000000000000;
        	9'b1_0000_0010:  	OUT <= 32'b11111100000000000000000000000000;

        	9'b1_0001_0011:  	OUT <= 32'b00000011000000000000000000000000;
        	9'b1_0010_0011:  	OUT <= 32'b00001111000000000000000000000000;
        	9'b1_0011_0011:  	OUT <= 32'b00111111000000000000000000000000;
        	9'b1_0100_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_0101_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_0110_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_0111_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1000_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1001_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1010_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1011_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1100_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1101_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1110_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_1111_0011:  	OUT <= 32'b11111111000000000000000000000000;
        	9'b1_0000_0011:  	OUT <= 32'b11111111000000000000000000000000;

        	9'b1_0001_0100:  	OUT <= 32'b00000000110000000000000000000000;
        	9'b1_0010_0100:  	OUT <= 32'b00000011110000000000000000000000;
        	9'b1_0011_0100:  	OUT <= 32'b00001111110000000000000000000000;
        	9'b1_0100_0100:  	OUT <= 32'b00111111110000000000000000000000;
        	9'b1_0101_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_0110_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_0111_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1000_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1001_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1010_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1011_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1100_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1101_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1110_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_1111_0100:  	OUT <= 32'b11111111110000000000000000000000;
        	9'b1_0000_0100:  	OUT <= 32'b11111111110000000000000000000000;

        	9'b1_0001_0101:  	OUT <= 32'b00000000001100000000000000000000;
        	9'b1_0010_0101:  	OUT <= 32'b00000000111100000000000000000000;
        	9'b1_0011_0101:  	OUT <= 32'b00000011111100000000000000000000;
        	9'b1_0100_0101:  	OUT <= 32'b00001111111100000000000000000000;
        	9'b1_0101_0101:  	OUT <= 32'b00111111111100000000000000000000;
        	9'b1_0110_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_0111_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1000_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1001_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1010_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1011_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1100_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1101_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1110_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_1111_0101:  	OUT <= 32'b11111111111100000000000000000000;
        	9'b1_0000_0101:  	OUT <= 32'b11111111111100000000000000000000;

        	9'b1_0001_0110:  	OUT <= 32'b00000000000011000000000000000000;
        	9'b1_0010_0110:  	OUT <= 32'b00000000001111000000000000000000;
        	9'b1_0011_0110:  	OUT <= 32'b00000000111111000000000000000000;
        	9'b1_0100_0110:  	OUT <= 32'b00000011111111000000000000000000;
        	9'b1_0101_0110:  	OUT <= 32'b00001111111111000000000000000000;
        	9'b1_0110_0110:  	OUT <= 32'b00111111111111000000000000000000;
        	9'b1_0111_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1000_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1001_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1010_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1011_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1100_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1101_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1110_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_1111_0110:  	OUT <= 32'b11111111111111000000000000000000;
        	9'b1_0000_0110:  	OUT <= 32'b11111111111111000000000000000000;

        	9'b1_0001_0111:  	OUT <= 32'b00000000000000110000000000000000;
        	9'b1_0010_0111:  	OUT <= 32'b00000000000011110000000000000000;
        	9'b1_0011_0111:  	OUT <= 32'b00000000001111110000000000000000;
        	9'b1_0100_0111:  	OUT <= 32'b00000000111111110000000000000000;
        	9'b1_0101_0111:  	OUT <= 32'b00000011111111110000000000000000;
        	9'b1_0110_0111:  	OUT <= 32'b00001111111111110000000000000000;
        	9'b1_0111_0111:  	OUT <= 32'b00111111111111110000000000000000;
        	9'b1_1000_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1001_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1010_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1011_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1100_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1101_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1110_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_1111_0111:  	OUT <= 32'b11111111111111110000000000000000;
        	9'b1_0000_0111:  	OUT <= 32'b11111111111111110000000000000000;

        	9'b1_0001_1000:  	OUT <= 32'b00000000000000001100000000000000;
        	9'b1_0010_1000:  	OUT <= 32'b00000000000000111100000000000000;
        	9'b1_0011_1000:  	OUT <= 32'b00000000000011111100000000000000;
        	9'b1_0100_1000:  	OUT <= 32'b00000000001111111100000000000000;
        	9'b1_0101_1000:  	OUT <= 32'b00000000111111111100000000000000;
        	9'b1_0110_1000:  	OUT <= 32'b00000011111111111100000000000000;
        	9'b1_0111_1000:  	OUT <= 32'b00001111111111111100000000000000;
        	9'b1_1000_1000:  	OUT <= 32'b00111111111111111100000000000000;
        	9'b1_1001_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1010_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1011_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1100_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1101_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1110_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_1111_1000:  	OUT <= 32'b11111111111111111100000000000000;
        	9'b1_0000_1000:  	OUT <= 32'b11111111111111111100000000000000;

        	9'b1_0001_1001:  	OUT <= 32'b00000000000000000011000000000000;
        	9'b1_0010_1001:  	OUT <= 32'b00000000000000001111000000000000;
        	9'b1_0011_1001:  	OUT <= 32'b00000000000000111111000000000000;
        	9'b1_0100_1001:  	OUT <= 32'b00000000000011111111000000000000;
        	9'b1_0101_1001:  	OUT <= 32'b00000000001111111111000000000000;
        	9'b1_0110_1001:  	OUT <= 32'b00000000111111111111000000000000;
        	9'b1_0111_1001:  	OUT <= 32'b00000011111111111111000000000000;
        	9'b1_1000_1001:  	OUT <= 32'b00001111111111111111000000000000;
        	9'b1_1001_1001:  	OUT <= 32'b00111111111111111111000000000000;
        	9'b1_1010_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_1011_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_1100_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_1101_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_1110_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_1111_1001:  	OUT <= 32'b11111111111111111111000000000000;
        	9'b1_0000_1001:  	OUT <= 32'b11111111111111111111000000000000;

        	9'b1_0001_1010:  	OUT <= 32'b00000000000000000000110000000000;
        	9'b1_0010_1010:  	OUT <= 32'b00000000000000000011110000000000;
        	9'b1_0011_1010:  	OUT <= 32'b00000000000000001111110000000000;
        	9'b1_0100_1010:  	OUT <= 32'b00000000000000111111110000000000;
        	9'b1_0101_1010:  	OUT <= 32'b00000000000011111111110000000000;
        	9'b1_0110_1010:  	OUT <= 32'b00000000001111111111110000000000;
        	9'b1_0111_1010:  	OUT <= 32'b00000000111111111111110000000000;
        	9'b1_1000_1010:  	OUT <= 32'b00000011111111111111110000000000;
        	9'b1_1001_1010:  	OUT <= 32'b00001111111111111111110000000000;
        	9'b1_1010_1010:  	OUT <= 32'b00111111111111111111110000000000;
        	9'b1_1011_1010:  	OUT <= 32'b11111111111111111111110000000000;
        	9'b1_1100_1010:  	OUT <= 32'b11111111111111111111110000000000;
        	9'b1_1101_1010:  	OUT <= 32'b11111111111111111111110000000000;
        	9'b1_1110_1010:  	OUT <= 32'b11111111111111111111110000000000;
        	9'b1_1111_1010:  	OUT <= 32'b11111111111111111111110000000000;
        	9'b1_0000_1010:  	OUT <= 32'b11111111111111111111110000000000;

        	9'b1_0001_1011:  	OUT <= 32'b00000000000000000000001100000000;
        	9'b1_0010_1011:  	OUT <= 32'b00000000000000000000111100000000;
        	9'b1_0011_1011:  	OUT <= 32'b00000000000000000011111100000000;
        	9'b1_0100_1011:  	OUT <= 32'b00000000000000001111111100000000;
        	9'b1_0101_1011:  	OUT <= 32'b00000000000000111111111100000000;
        	9'b1_0110_1011:  	OUT <= 32'b00000000000011111111111100000000;
        	9'b1_0111_1011:  	OUT <= 32'b00000000001111111111111100000000;
        	9'b1_1000_1011:  	OUT <= 32'b00000000111111111111111100000000;
        	9'b1_1001_1011:  	OUT <= 32'b00000011111111111111111100000000;
        	9'b1_1010_1011:  	OUT <= 32'b00001111111111111111111100000000;
        	9'b1_1011_1011:  	OUT <= 32'b00111111111111111111111100000000;
        	9'b1_1100_1011:  	OUT <= 32'b11111111111111111111111100000000;
        	9'b1_1101_1011:  	OUT <= 32'b11111111111111111111111100000000;
        	9'b1_1110_1011:  	OUT <= 32'b11111111111111111111111100000000;
        	9'b1_1111_1011:  	OUT <= 32'b11111111111111111111111100000000;
        	9'b1_0000_1011:  	OUT <= 32'b11111111111111111111111100000000;

        	9'b1_0001_1100:  	OUT <= 32'b00000000000000000000000011000000;
        	9'b1_0010_1100:  	OUT <= 32'b00000000000000000000001111000000;
        	9'b1_0011_1100:  	OUT <= 32'b00000000000000000000111111000000;
        	9'b1_0100_1100:  	OUT <= 32'b00000000000000000011111111000000;
        	9'b1_0101_1100:  	OUT <= 32'b00000000000000001111111111000000;
        	9'b1_0110_1100:  	OUT <= 32'b00000000000000111111111111000000;
        	9'b1_0111_1100:  	OUT <= 32'b00000000000011111111111111000000;
        	9'b1_1000_1100:  	OUT <= 32'b00000000001111111111111111000000;
        	9'b1_1001_1100:  	OUT <= 32'b00000000111111111111111111000000;
        	9'b1_1010_1100:  	OUT <= 32'b00000011111111111111111111000000;
        	9'b1_1011_1100:  	OUT <= 32'b00001111111111111111111111000000;
        	9'b1_1100_1100:  	OUT <= 32'b00111111111111111111111111000000;
        	9'b1_1101_1100:  	OUT <= 32'b11111111111111111111111111000000;
        	9'b1_1110_1100:  	OUT <= 32'b11111111111111111111111111000000;
        	9'b1_1111_1100:  	OUT <= 32'b11111111111111111111111111000000;
        	9'b1_0000_1100:  	OUT <= 32'b11111111111111111111111111000000;

        	9'b1_0001_1101:  	OUT <= 32'b00000000000000000000000000110000;
        	9'b1_0010_1101:  	OUT <= 32'b00000000000000000000000011110000;
        	9'b1_0011_1101:  	OUT <= 32'b00000000000000000000001111110000;
        	9'b1_0100_1101:  	OUT <= 32'b00000000000000000000111111110000;
        	9'b1_0101_1101:  	OUT <= 32'b00000000000000000011111111110000;
        	9'b1_0110_1101:  	OUT <= 32'b00000000000000001111111111110000;
        	9'b1_0111_1101:  	OUT <= 32'b00000000000000111111111111110000;
        	9'b1_1000_1101:  	OUT <= 32'b00000000000011111111111111110000;
        	9'b1_1001_1101:  	OUT <= 32'b00000000001111111111111111110000;
        	9'b1_1010_1101:  	OUT <= 32'b00000000111111111111111111110000;
        	9'b1_1011_1101:  	OUT <= 32'b00000011111111111111111111110000;
        	9'b1_1100_1101:  	OUT <= 32'b00001111111111111111111111110000;
        	9'b1_1101_1101:  	OUT <= 32'b00111111111111111111111111110000;
        	9'b1_1110_1101:  	OUT <= 32'b11111111111111111111111111110000;
        	9'b1_1111_1101:  	OUT <= 32'b11111111111111111111111111110000;
        	9'b1_0000_1101:  	OUT <= 32'b11111111111111111111111111110000;

        	9'b1_0001_1110:  	OUT <= 32'b00000000000000000000000000001100;
        	9'b1_0010_1110:  	OUT <= 32'b00000000000000000000000000111100;
        	9'b1_0011_1110:  	OUT <= 32'b00000000000000000000000011111100;
        	9'b1_0100_1110:  	OUT <= 32'b00000000000000000000001111111100;
        	9'b1_0101_1110:  	OUT <= 32'b00000000000000000000111111111100;
        	9'b1_0110_1110:  	OUT <= 32'b00000000000000000011111111111100;
        	9'b1_0111_1110:  	OUT <= 32'b00000000000000001111111111111100;
        	9'b1_1000_1110:  	OUT <= 32'b00000000000000111111111111111100;
        	9'b1_1001_1110:  	OUT <= 32'b00000000000011111111111111111100;
        	9'b1_1010_1110:  	OUT <= 32'b00000000001111111111111111111100;
        	9'b1_1011_1110:  	OUT <= 32'b00000000111111111111111111111100;
        	9'b1_1100_1110:  	OUT <= 32'b00000011111111111111111111111100;
        	9'b1_1101_1110:  	OUT <= 32'b00001111111111111111111111111100;
        	9'b1_1110_1110:  	OUT <= 32'b00111111111111111111111111111100;
        	9'b1_1111_1110:  	OUT <= 32'b11111111111111111111111111111100;
        	9'b1_0000_1110:  	OUT <= 32'b11111111111111111111111111111100;

        	9'b1_0001_1111:  	OUT <= 32'b00000000000000000000000000000011;
        	9'b1_0010_1111:  	OUT <= 32'b00000000000000000000000000001111;
        	9'b1_0011_1111:  	OUT <= 32'b00000000000000000000000000111111;
        	9'b1_0100_1111:  	OUT <= 32'b00000000000000000000000011111111;
        	9'b1_0101_1111:  	OUT <= 32'b00000000000000000000001111111111;
        	9'b1_0110_1111:  	OUT <= 32'b00000000000000000000111111111111;
        	9'b1_0111_1111:  	OUT <= 32'b00000000000000000011111111111111;
        	9'b1_1000_1111:  	OUT <= 32'b00000000000000001111111111111111;
        	9'b1_1001_1111:  	OUT <= 32'b00000000000000111111111111111111;
        	9'b1_1010_1111:  	OUT <= 32'b00000000000011111111111111111111;
        	9'b1_1011_1111:  	OUT <= 32'b00000000001111111111111111111111;
        	9'b1_1100_1111:  	OUT <= 32'b00000000111111111111111111111111;
        	9'b1_1101_1111:  	OUT <= 32'b00000011111111111111111111111111;
        	9'b1_1110_1111:  	OUT <= 32'b00001111111111111111111111111111;
        	9'b1_1111_1111:  	OUT <= 32'b00111111111111111111111111111111;
        	9'b1_0000_1111:  	OUT <= 32'b11111111111111111111111111111111;
        endcase
    end
endmodule

/***************************************************************
 * 4BPP テーブル
 ***************************************************************/
module T9990_BLIT_BITMASK_4BPP (
    input wire          CLK,
    input wire          DIX,
    input wire [2:0]    OFFSET,
    input wire [2:0]    COUNT,
    output reg [31:0]   OUT
)/* synthesis syn_romstyle="block_rom" */;
    always_ff @(posedge CLK) begin
        case ({DIX,COUNT[2:0],OFFSET[2:0]})
        	7'b0_001_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b0_010_000:       OUT <= 32'b11111111000000000000000000000000;
        	7'b0_011_000:       OUT <= 32'b11111111111100000000000000000000;
        	7'b0_100_000:       OUT <= 32'b11111111111111110000000000000000;
        	7'b0_101_000:       OUT <= 32'b11111111111111111111000000000000;
        	7'b0_110_000:       OUT <= 32'b11111111111111111111111100000000;
        	7'b0_111_000:       OUT <= 32'b11111111111111111111111111110000;
        	7'b0_000_000:       OUT <= 32'b11111111111111111111111111111111;

        	7'b0_001_001:       OUT <= 32'b00001111000000000000000000000000;
        	7'b0_010_001:       OUT <= 32'b00001111111100000000000000000000;
        	7'b0_011_001:       OUT <= 32'b00001111111111110000000000000000;
        	7'b0_100_001:       OUT <= 32'b00001111111111111111000000000000;
        	7'b0_101_001:       OUT <= 32'b00001111111111111111111100000000;
        	7'b0_110_001:       OUT <= 32'b00001111111111111111111111110000;
        	7'b0_111_001:       OUT <= 32'b00001111111111111111111111111111;
        	7'b0_000_001:       OUT <= 32'b00001111111111111111111111111111;

        	7'b0_001_010:       OUT <= 32'b00000000111100000000000000000000;
        	7'b0_010_010:       OUT <= 32'b00000000111111110000000000000000;
        	7'b0_011_010:       OUT <= 32'b00000000111111111111000000000000;
        	7'b0_100_010:       OUT <= 32'b00000000111111111111111100000000;
        	7'b0_101_010:       OUT <= 32'b00000000111111111111111111110000;
        	7'b0_110_010:       OUT <= 32'b00000000111111111111111111111111;
        	7'b0_111_010:       OUT <= 32'b00000000111111111111111111111111;
        	7'b0_000_010:       OUT <= 32'b00000000111111111111111111111111;

        	7'b0_001_011:       OUT <= 32'b00000000000011110000000000000000;
        	7'b0_010_011:       OUT <= 32'b00000000000011111111000000000000;
        	7'b0_011_011:       OUT <= 32'b00000000000011111111111100000000;
        	7'b0_100_011:       OUT <= 32'b00000000000011111111111111110000;
        	7'b0_101_011:       OUT <= 32'b00000000000011111111111111111111;
        	7'b0_110_011:       OUT <= 32'b00000000000011111111111111111111;
        	7'b0_111_011:       OUT <= 32'b00000000000011111111111111111111;
        	7'b0_000_011:       OUT <= 32'b00000000000011111111111111111111;

        	7'b0_001_100:       OUT <= 32'b00000000000000001111000000000000;
        	7'b0_010_100:       OUT <= 32'b00000000000000001111111100000000;
        	7'b0_011_100:       OUT <= 32'b00000000000000001111111111110000;
        	7'b0_100_100:       OUT <= 32'b00000000000000001111111111111111;
        	7'b0_101_100:       OUT <= 32'b00000000000000001111111111111111;
        	7'b0_110_100:       OUT <= 32'b00000000000000001111111111111111;
        	7'b0_111_100:       OUT <= 32'b00000000000000001111111111111111;
        	7'b0_000_100:       OUT <= 32'b00000000000000001111111111111111;

        	7'b0_001_101:       OUT <= 32'b00000000000000000000111100000000;
        	7'b0_010_101:       OUT <= 32'b00000000000000000000111111110000;
        	7'b0_011_101:       OUT <= 32'b00000000000000000000111111111111;
        	7'b0_100_101:       OUT <= 32'b00000000000000000000111111111111;
        	7'b0_101_101:       OUT <= 32'b00000000000000000000111111111111;
        	7'b0_110_101:       OUT <= 32'b00000000000000000000111111111111;
        	7'b0_111_101:       OUT <= 32'b00000000000000000000111111111111;
        	7'b0_000_101:       OUT <= 32'b00000000000000000000111111111111;

        	7'b0_001_110:       OUT <= 32'b00000000000000000000000011110000;
        	7'b0_010_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_011_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_100_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_101_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_110_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_111_110:       OUT <= 32'b00000000000000000000000011111111;
        	7'b0_000_110:       OUT <= 32'b00000000000000000000000011111111;

        	7'b0_001_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_010_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_011_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_100_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_101_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_110_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_111_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b0_000_111:       OUT <= 32'b00000000000000000000000000001111;

        	7'b1_001_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_010_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_011_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_100_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_101_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_110_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_111_000:       OUT <= 32'b11110000000000000000000000000000;
        	7'b1_000_000:       OUT <= 32'b11110000000000000000000000000000;

        	7'b1_001_001:       OUT <= 32'b00001111000000000000000000000000;
        	7'b1_010_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_011_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_100_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_101_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_110_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_111_001:       OUT <= 32'b11111111000000000000000000000000;
        	7'b1_000_001:       OUT <= 32'b11111111000000000000000000000000;

        	7'b1_001_010:       OUT <= 32'b00000000111100000000000000000000;
        	7'b1_010_010:       OUT <= 32'b00001111111100000000000000000000;
        	7'b1_011_010:       OUT <= 32'b11111111111100000000000000000000;
        	7'b1_100_010:       OUT <= 32'b11111111111100000000000000000000;
        	7'b1_101_010:       OUT <= 32'b11111111111100000000000000000000;
        	7'b1_110_010:       OUT <= 32'b11111111111100000000000000000000;
        	7'b1_111_010:       OUT <= 32'b11111111111100000000000000000000;
        	7'b1_000_010:       OUT <= 32'b11111111111100000000000000000000;

        	7'b1_001_011:       OUT <= 32'b00000000000011110000000000000000;
        	7'b1_010_011:       OUT <= 32'b00000000111111110000000000000000;
        	7'b1_011_011:       OUT <= 32'b00001111111111110000000000000000;
        	7'b1_100_011:       OUT <= 32'b11111111111111110000000000000000;
        	7'b1_101_011:       OUT <= 32'b11111111111111110000000000000000;
        	7'b1_110_011:       OUT <= 32'b11111111111111110000000000000000;
        	7'b1_111_011:       OUT <= 32'b11111111111111110000000000000000;
        	7'b1_000_011:       OUT <= 32'b11111111111111110000000000000000;

        	7'b1_001_100:       OUT <= 32'b00000000000000001111000000000000;
        	7'b1_010_100:       OUT <= 32'b00000000000011111111000000000000;
        	7'b1_011_100:       OUT <= 32'b00000000111111111111000000000000;
        	7'b1_100_100:       OUT <= 32'b00001111111111111111000000000000;
        	7'b1_101_100:       OUT <= 32'b11111111111111111111000000000000;
        	7'b1_110_100:       OUT <= 32'b11111111111111111111000000000000;
        	7'b1_111_100:       OUT <= 32'b11111111111111111111000000000000;
        	7'b1_000_100:       OUT <= 32'b11111111111111111111000000000000;

        	7'b1_001_101:       OUT <= 32'b00000000000000000000111100000000;
        	7'b1_010_101:       OUT <= 32'b00000000000000001111111100000000;
        	7'b1_011_101:       OUT <= 32'b00000000000011111111111100000000;
        	7'b1_100_101:       OUT <= 32'b00000000111111111111111100000000;
        	7'b1_101_101:       OUT <= 32'b00001111111111111111111100000000;
        	7'b1_110_101:       OUT <= 32'b11111111111111111111111100000000;
        	7'b1_111_101:       OUT <= 32'b11111111111111111111111100000000;
        	7'b1_000_101:       OUT <= 32'b11111111111111111111111100000000;

        	7'b1_001_110:       OUT <= 32'b00000000000000000000000011110000;
        	7'b1_010_110:       OUT <= 32'b00000000000000000000111111110000;
        	7'b1_011_110:       OUT <= 32'b00000000000000001111111111110000;
        	7'b1_100_110:       OUT <= 32'b00000000000011111111111111110000;
        	7'b1_101_110:       OUT <= 32'b00000000111111111111111111110000;
        	7'b1_110_110:       OUT <= 32'b00001111111111111111111111110000;
        	7'b1_111_110:       OUT <= 32'b11111111111111111111111111110000;
        	7'b1_000_110:       OUT <= 32'b11111111111111111111111111110000;

        	7'b1_001_111:       OUT <= 32'b00000000000000000000000000001111;
        	7'b1_010_111:       OUT <= 32'b00000000000000000000000011111111;
        	7'b1_011_111:       OUT <= 32'b00000000000000000000111111111111;
        	7'b1_100_111:       OUT <= 32'b00000000000000001111111111111111;
        	7'b1_101_111:       OUT <= 32'b00000000000011111111111111111111;
        	7'b1_110_111:       OUT <= 32'b00000000111111111111111111111111;
        	7'b1_111_111:       OUT <= 32'b00001111111111111111111111111111;
        	7'b1_000_111:       OUT <= 32'b11111111111111111111111111111111;
        endcase
    end
endmodule

/***************************************************************
 * 8BPP テーブル
 ***************************************************************/
module T9990_BLIT_BITMASK_8BPP (
    input wire          CLK,
    input wire          DIX,
    input wire [1:0]    OFFSET,
    input wire [1:0]    COUNT,
    output reg [31:0]   OUT
)/* synthesis syn_romstyle="block_rom" */;
    always_ff @(posedge CLK) begin
        case ({DIX,COUNT[1:0],OFFSET[1:0]})
        	5'b0_01_00:         OUT <= 32'b11111111000000000000000000000000;
        	5'b0_10_00:         OUT <= 32'b11111111111111110000000000000000;
        	5'b0_11_00:         OUT <= 32'b11111111111111111111111100000000;
        	5'b0_00_00:         OUT <= 32'b11111111111111111111111111111111;

        	5'b0_01_01:         OUT <= 32'b00000000111111110000000000000000;
        	5'b0_10_01:         OUT <= 32'b00000000111111111111111100000000;
        	5'b0_11_01:         OUT <= 32'b00000000111111111111111111111111;
        	5'b0_00_01:         OUT <= 32'b00000000111111111111111111111111;

        	5'b0_01_10:         OUT <= 32'b00000000000000001111111100000000;
        	5'b0_10_10:         OUT <= 32'b00000000000000001111111111111111;
        	5'b0_11_10:         OUT <= 32'b00000000000000001111111111111111;
        	5'b0_00_10:         OUT <= 32'b00000000000000001111111111111111;

        	5'b0_01_11:         OUT <= 32'b00000000000000000000000011111111;
        	5'b0_10_11:         OUT <= 32'b00000000000000000000000011111111;
        	5'b0_11_11:         OUT <= 32'b00000000000000000000000011111111;
        	5'b0_00_11:         OUT <= 32'b00000000000000000000000011111111;

        	5'b1_01_00:         OUT <= 32'b11111111000000000000000000000000;
        	5'b1_10_00:         OUT <= 32'b11111111000000000000000000000000;
        	5'b1_11_00:         OUT <= 32'b11111111000000000000000000000000;
        	5'b1_00_00:         OUT <= 32'b11111111000000000000000000000000;

        	5'b1_01_01:         OUT <= 32'b00000000111111110000000000000000;
        	5'b1_10_01:         OUT <= 32'b11111111111111110000000000000000;
        	5'b1_11_01:         OUT <= 32'b11111111111111110000000000000000;
        	5'b1_00_01:         OUT <= 32'b11111111111111110000000000000000;

        	5'b1_01_10:         OUT <= 32'b00000000000000001111111100000000;
        	5'b1_10_10:         OUT <= 32'b00000000111111111111111100000000;
        	5'b1_11_10:         OUT <= 32'b11111111111111111111111100000000;
        	5'b1_00_10:         OUT <= 32'b11111111111111111111111100000000;

        	5'b1_01_11:         OUT <= 32'b00000000000000000000000011111111;
        	5'b1_10_11:         OUT <= 32'b00000000000000001111111111111111;
        	5'b1_11_11:         OUT <= 32'b00000000111111111111111111111111;
        	5'b1_00_11:         OUT <= 32'b11111111111111111111111111111111;
        endcase
    end
endmodule

/***************************************************************
 * 16BPP テーブル
 ***************************************************************/
module T9990_BLIT_BITMASK_16BPP (
    input wire          CLK,
    input wire          DIX,
    input wire [0:0]    OFFSET,
    input wire [0:0]    COUNT,
    output reg [31:0]   OUT
)/* synthesis syn_romstyle="block_rom" */;
    always_ff @(posedge CLK) begin
        case ({DIX,COUNT[0:0],OFFSET[0:0]})
        	3'b0_1_0:           OUT <= 32'b11111111111111110000000000000000;
        	3'b0_0_0:           OUT <= 32'b11111111111111111111111111111111;

        	3'b0_1_1:           OUT <= 32'b00000000000000001111111111111111;
        	3'b0_0_1:           OUT <= 32'b00000000000000001111111111111111;

        	3'b1_1_0:           OUT <= 32'b11111111111111110000000000000000;
        	3'b1_0_0:           OUT <= 32'b11111111111111110000000000000000;

        	3'b1_1_1:           OUT <= 32'b00000000000000001111111111111111;
        	3'b1_0_1:           OUT <= 32'b11111111111111111111111111111111;
        endcase
    end
endmodule

`default_nettype wire
